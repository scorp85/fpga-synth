module sample(index, clk, saida);
	input [2:0] index;
	input clk;
	output reg[7:0] saida;
endmodule

